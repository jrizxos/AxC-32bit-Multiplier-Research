signal s10060,s10059,s10058,s10057,s10056,s10055,s10054,s10053,s10052,--STAGE1
s10051,s10050,s10049,s10048,s10047,s10046,s10045,s10044,s10043,s10042,
s10041,s10040,s10039,s10038,s10037,s10036,s10035,s10034,s10033,s10032,
s10031,s10030,s10029,s10028,s10027,s10026,s10025,s10024,s10023,s10022,
s10021,s10020,s10019,s10018,s10017,s10016,s10015,s10014,s10013,s10012,
s10011,s10010,s10009,s10008,s10007,s10006,s10005,s10004,s10003,s10002,
s10157,s10156,s10155,s10154,s10153,s10152,s10151,s10150,s10149,s10148,
s10147,s10146,s10145,s10144,s10143,s10142,s10141,s10140,s10139,s10138,
s10137,s10136,s10135,s10134,s10133,s10132,s10131,s10130,s10129,s10128,
s10127,s10126,s10125,s10124,s10123,s10122,s10121,s10120,s10119,s10118,
s10117,s10116,s10115,s10114,s10113,s10112,s10111,s10110,s10109,s10108,
s10107,s10106,s10105,s10254,s10253,s10252,s10251,s10250,s10249,s10248,
s10247,s10246,s10245,s10244,s10243,s10242,s10241,s10240,s10239,s10238,
s10237,s10236,s10235,s10234,s10233,s10232,s10231,s10230,s10229,s10228,
s10227,s10226,s10225,s10224,s10223,s10222,s10221,s10220,s10219,s10218,
s10217,s10216,s10215,s10214,s10213,s10212,s10211,s10210,s10209,s10208,
s10351,s10350,s10349,s10348,s10347,s10346,s10345,s10344,s10343,s10342,
s10341,s10340,s10339,s10338,s10337,s10336,s10335,s10334,s10333,s10332,
s10331,s10330,s10329,s10328,s10327,s10326,s10325,s10324,s10323,s10322,
s10321,s10320,s10319,s10318,s10317,s10316,s10315,s10314,s10313,s10312,
s10311,s10448,s10447,s10446,s10445,s10444,s10443,s10442,s10441,s10440,
s10439,s10438,s10437,s10436,s10435,s10434,s10433,s10432,s10431,s10430,
s10429,s10428,s10427,s10426,s10425,s10424,s10423,s10422,s10421,s10420,
s10419,s10418,s10417,s10416,s10415,s10414,s10545,s10544,s10543,s10542,
s10541,s10540,s10539,s10538,s10537,s10536,s10535,s10534,s10533,s10532,
s10531,s10530,s10529,s10528,s10527,s10526,s10525,s10524,s10523,s10522,
s10521,s10520,s10519,s10518,s10517,s10642,s10641,s10640,s10639,s10638,
s10637,s10636,s10635,s10634,s10633,s10632,s10631,s10630,s10629,s10628,
s10627,s10626,s10625,s10624,s10623,s10622,s10621,s10620,s10739,s10738,
s10737,s10736,s10735,s10734,s10733,s10732,s10731,s10730,s10729,s10728,
s10727,s10726,s10725,s10724,s10723,s10836,s10835,s10834,s10833,s10832,
s10831,s10830,s10829,s10828,s10827,s10826,s10933,s10932,s10931,s10930,
s10929,

s20061,s20059,s20058,s20057,s20056,s20055,s20054,s20053,s20052,s20051,--STAGE2
s20050,s20049,s20048,s20047,s20046,s20045,s20044,s20043,s20042,s20041,
s20040,s20039,s20038,s20037,s20036,s20035,s20034,s20033,s20032,s20031,
s20030,s20029,s20028,s20027,s20026,s20025,s20024,s20023,s20022,s20021,
s20020,s20019,s20018,s20017,s20016,s20015,s20014,s20013,s20012,s20011,
s20010,s20009,s20008,s20007,s20006,s20005,s20004,s20003,s20155,s20154,
s20153,s20152,s20151,s20150,s20149,s20148,s20147,s20146,s20145,s20144,
s20143,s20142,s20141,s20140,s20139,s20138,s20137,s20136,s20135,s20134,
s20133,s20132,s20131,s20130,s20129,s20128,s20127,s20126,s20125,s20124,
s20123,s20122,s20121,s20120,s20119,s20118,s20117,s20116,s20115,s20114,
s20113,s20112,s20111,s20110,s20109,s20107,s20252,s20250,s20249,s20248,
s20247,s20246,s20245,s20244,s20243,s20242,s20241,s20240,s20239,s20238,
s20237,s20236,s20235,s20234,s20233,s20232,s20231,s20230,s20229,s20228,
s20227,s20226,s20225,s20224,s20223,s20222,s20221,s20220,s20219,s20218,
s20217,s20216,s20215,s20214,s20213,s20212,s20346,s20345,s20344,s20343,
s20342,s20341,s20340,s20339,s20338,s20337,s20336,s20335,s20334,s20333,
s20332,s20331,s20330,s20329,s20328,s20327,s20326,s20325,s20324,s20323,
s20322,s20321,s20320,s20319,s20318,s20316,s20443,s20441,s20440,s20439,
s20438,s20437,s20436,s20435,s20434,s20433,s20432,s20431,s20430,s20429,
s20428,s20427,s20426,s20425,s20424,s20423,s20422,s20421,s20537,s20536,
s20535,s20534,s20533,s20532,s20531,s20530,s20529,s20528,s20527,s20525,
s20634,s20632,s20631,s20630,

s30060,s30059,s30058,s30057,s30056,s30055,s30054,s30053,s30052,s30051,--STAGE3
s30050,s30049,s30048,s30047,s30046,s30045,s30044,s30043,s30042,s30041,
s30040,s30039,s30038,s30037,s30036,s30035,s30034,s30033,s30032,s30031,
s30030,s30029,s30028,s30027,s30026,s30025,s30024,s30023,s30022,s30021,
s30020,s30019,s30018,s30017,s30016,s30015,s30014,s30013,s30012,s30011,
s30010,s30009,s30008,s30007,s30006,s30005,s30004,s30156,s30155,s30153,
s30152,s30151,s30150,s30149,s30148,s30147,s30146,s30145,s30144,s30143,
s30142,s30141,s30140,s30139,s30138,s30137,s30136,s30135,s30134,s30133,
s30132,s30131,s30130,s30129,s30128,s30127,s30126,s30125,s30124,s30123,
s30122,s30121,s30120,s30119,s30118,s30117,s30116,s30115,s30114,s30113,
s30112,s30111,s30110,s30108,s30249,s30247,s30246,s30245,s30244,s30243,
s30242,s30241,s30240,s30239,s30238,s30237,s30236,s30235,s30234,s30233,
s30232,s30231,s30230,s30229,s30228,s30227,s30226,s30225,s30224,s30223,
s30222,s30221,s30220,s30219,s30218,s30217,s30215,s30342,s30340,s30339,
s30338,s30337,s30336,s30335,s30334,s30333,s30332,s30331,s30330,s30329,
s30328,s30327,s30326,s30325,s30324,s30322,s30435,s30433,s30432,s30431,
s30428,

s40058,s40057,s40056,s40055,s40054,s40053,s40052,s40051,s40050,s40049,--STAGE4
s40048,s40047,s40046,s40045,s40044,s40043,s40042,s40041,s40040,s40039,
s40038,s40037,s40036,s40035,s40034,s40033,s40032,s40031,s40030,s40029,
s40028,s40027,s40026,s40025,s40024,s40023,s40022,s40021,s40020,s40019,
s40018,s40017,s40016,s40015,s40014,s40013,s40012,s40011,s40010,s40009,
s40008,s40006,s40148,s40147,s40146,s40145,s40144,s40143,s40142,s40141,
s40140,s40139,s40138,s40137,s40136,s40135,s40134,s40133,s40132,s40131,
s40130,s40129,s40128,s40127,s40126,s40125,s40124,s40123,s40122,s40121,
s40120,s40119,s40118,s40116,s40238,s40237,s40236,s40235,s40234,s40233,
s40232,s40231,s40230,s40229,s40228,s40226,

s50059,s50056,s50054,s50053,s50052,s50051,s50050,s50049,s50048,s50047,--STAGE5
s50046,s50045,s50044,s50043,s50042,s50041,s50040,s50039,s50038,s50037,
s50036,s50035,s50034,s50033,s50032,s50031,s50030,s50029,s50028,s50027,
s50026,s50025,s50024,s50023,s50022,s50021,s50020,s50019,s50018,s50017,
s50016,s50015,s50014,s50013,s50012,s50011,s50009,s50007,s50141,s50140,
s50139,s50138,s50137,s50136,s50135,s50134,s50133,s50132,s50131,s50130,
s50129,s50127,s50125,s50123,

s60060,s60057,s60055,s60051,s60050,s60049,s60048,s60047,s60046,s60045,--STAGE6
s60044,s60043,s60042,s60041,s60040,s60039,s60038,s60037,s60036,s60035,
s60034,s60033,s60032,s60031,s60030,s60029,s60028,s60027,s60026,s60025,
s60024,s60023,s60022,s60021,s60020,s60019,s60017,s60015,s60013,s60010,

s70061,s70058,s70052,s70049,s70044,s70043,s70042,s70041,s70040,s70039,--STAGE7
s70038,s70037,s70036,s70035,s70034,s70033,s70032,s70031,s70030,s70029,
s70028,s70027,s70026,s70024,s70022,s70018,s70016,s70014,

s80062,s80054,s80053,s80051,s80050,s80048,s80047,s80046,s80045,s80044,--STAGE8
s80043,s80042,s80041,s80040,s80039,s80038,s80037,s80036,s80035,s80034,
s80033,s80032,s80031,s80030,s80029,s80028,s80027,s80026,s80025,s80024,
s80023,s80021,s80020,s80019,s80017												: std_logic; 

prodA(0)  <= p(0);
prodA(1)  <= p(1);
prodA(2)  <= s10002;
prodA(3)  <= s20003;
prodA(4)  <= s30004;
prodA(5)  <= s30005;
prodA(6)  <= s40006;
prodA(7)  <= s50007;
prodA(8)  <= s40008;
prodA(9)  <= s50009;
prodA(10) <= s60010;
prodA(11) <= s50011;
prodA(12) <= s50012;
prodA(13) <= s60013;
prodA(14) <= s70014;
prodA(15) <= s60015;
prodA(16) <= s70016;
prodA(17) <= s80017;
prodA(18) <= s70018;
prodA(19) <= s80019;
prodA(20) <= s80020;
prodA(21) <= s80021;
prodA(22) <= s70022;
prodA(23) <= s80023;
prodA(24) <= s80024;
prodA(25) <= s80025;
prodA(26) <= s80026;
prodA(27) <= s80027;
prodA(28) <= s80028;
prodA(29) <= s80029;
prodA(30) <= s80030;
prodA(31) <= s80031;
prodA(32) <= s80032;
prodA(33) <= s80033;
prodA(34) <= s80034;
prodA(35) <= s80035;
prodA(36) <= s80036;
prodA(37) <= s80037;
prodA(38) <= s80038;
prodA(39) <= s80039;
prodA(40) <= s80040;
prodA(41) <= s80041;
prodA(42) <= s80042;
prodA(43) <= s80043;
prodA(44) <= s80044;
prodA(45) <= s80045;
prodA(46) <= s80046;
prodA(47) <= s80047;
prodA(48) <= s80048;
prodA(49) <= s70049;
prodA(50) <= s80050;
prodA(51) <= s80051;
prodA(52) <= s70052;
prodA(53) <= s80053;
prodA(54) <= s80054;
prodA(55) <= s60055;
prodA(56) <= s50056;
prodA(57) <= s60057;
prodA(58) <= s70058;
prodA(59) <= s50059;
prodA(60) <= s60060;
prodA(61) <= s70061;
prodA(62) <= s80062;
prodA(63) <= '0';

prodB(0)  <= '0';
prodB(1)  <= p(32);
prodB(2)  <= '0';
prodB(3)  <= '0';
prodB(4)  <= '0';
prodB(5)  <= c30004;
prodB(6)  <= '0';
prodB(7)  <= '0';
prodB(8)  <= c50007;
prodB(9)  <= '0';
prodB(10) <= '0';
prodB(11) <= c60010;
prodB(12) <= c50011;
prodB(13) <= '0';
prodB(14) <= '0';
prodB(15) <= c70014;
prodB(16) <= '0';
prodB(17) <= '0';
prodB(18) <= c80017;
prodB(19) <= '0';
prodB(20) <= c80019;
prodB(21) <= c80020;
prodB(22) <= c80021;
prodB(23) <= '0';
prodB(24) <= c80023;
prodB(25) <= c80024;
prodB(26) <= c80025;
prodB(27) <= c80026;
prodB(28) <= c80027;
prodB(29) <= c80028;
prodB(30) <= c80029;
prodB(31) <= c80030;
prodB(32) <= c80031;
prodB(33) <= c80032;
prodB(34) <= c80033;
prodB(35) <= c80034;
prodB(36) <= c80035;
prodB(37) <= c80036;
prodB(38) <= c80037;
prodB(39) <= c80038;
prodB(40) <= c80039;
prodB(41) <= c80040;
prodB(42) <= c80041;
prodB(43) <= c80042;
prodB(44) <= c80043;
prodB(45) <= c80044;
prodB(46) <= c80045;
prodB(47) <= c80046;
prodB(48) <= c80047;
prodB(49) <= c80048;
prodB(50) <= '0';
prodB(51) <= c80050;
prodB(52) <= c80051;
prodB(53) <= '0';
prodB(54) <= c80053;
prodB(55) <= c80054;
prodB(56) <= c60055;
prodB(57) <= '0';
prodB(58) <= '0';
prodB(59) <= c70058;
prodB(60) <= '0';
prodB(61) <= '0';
prodB(62) <= '0';
prodB(63) <= c80062;

--STAGE 1 -  FULL ADDERS:320 | HALF ADDERS:0
--GROUP 00
fa10002 : full_adder port map(p(2),p(33),p(64),s10002,c10002);
fa10003 : full_adder port map(p(3),p(34),p(65),s10003,c10003);
fa10004 : full_adder port map(p(4),p(35),p(66),s10004,c10004);
fa10005 : full_adder port map(p(5),p(36),p(67),s10005,c10005);
fa10006 : full_adder port map(p(6),p(37),p(68),s10006,c10006);
fa10007 : full_adder port map(p(7),p(38),p(69),s10007,c10007);
fa10008 : full_adder port map(p(8),p(39),p(70),s10008,c10008);
fa10009 : full_adder port map(p(9),p(40),p(71),s10009,c10009);
fa10010 : full_adder port map(p(10),p(41),p(72),s10010,c10010);
fa10011 : full_adder port map(p(11),p(42),p(73),s10011,c10011);
fa10012 : full_adder port map(p(12),p(43),p(74),s10012,c10012);
fa10013 : full_adder port map(p(13),p(44),p(75),s10013,c10013);
fa10014 : full_adder port map(p(14),p(45),p(76),s10014,c10014);
fa10015 : full_adder port map(p(15),p(46),p(77),s10015,c10015);
fa10016 : full_adder port map(p(16),p(47),p(78),s10016,c10016);
fa10017 : full_adder port map(p(17),p(48),p(79),s10017,c10017);
fa10018 : full_adder port map(p(18),p(49),p(80),s10018,c10018);
fa10019 : full_adder port map(p(19),p(50),p(81),s10019,c10019);
fa10020 : full_adder port map(p(20),p(51),p(82),s10020,c10020);
fa10021 : full_adder port map(p(21),p(52),p(83),s10021,c10021);
fa10022 : full_adder port map(p(22),p(53),p(84),s10022,c10022);
fa10023 : full_adder port map(p(23),p(54),p(85),s10023,c10023);
fa10024 : full_adder port map(p(24),p(55),p(86),s10024,c10024);
fa10025 : full_adder port map(p(25),p(56),p(87),s10025,c10025);
fa10026 : full_adder port map(p(26),p(57),p(88),s10026,c10026);
fa10027 : full_adder port map(p(27),p(58),p(89),s10027,c10027);
fa10028 : full_adder port map(p(28),p(59),p(90),s10028,c10028);
fa10029 : full_adder port map(p(29),p(60),p(91),s10029,c10029);
fa10030 : full_adder port map(p(30),p(61),p(92),s10030,c10030);
fa10031 : full_adder port map(p(31),p(62),p(93),s10031,c10031);
fa10032 : full_adder port map(p(63),p(94),p(125),s10032,c10032);
fa10033 : full_adder port map(p(95),p(126),p(157),s10033,c10033);
fa10034 : full_adder port map(p(127),p(158),p(189),s10034,c10034);
fa10035 : full_adder port map(p(159),p(190),p(221),s10035,c10035);
fa10036 : full_adder port map(p(191),p(222),p(253),s10036,c10036);
fa10037 : full_adder port map(p(223),p(254),p(285),s10037,c10037);
fa10038 : full_adder port map(p(255),p(286),p(317),s10038,c10038);
fa10039 : full_adder port map(p(287),p(318),p(349),s10039,c10039);
fa10040 : full_adder port map(p(319),p(350),p(381),s10040,c10040);
fa10041 : full_adder port map(p(351),p(382),p(413),s10041,c10041);
fa10042 : full_adder port map(p(383),p(414),p(445),s10042,c10042);
fa10043 : full_adder port map(p(415),p(446),p(477),s10043,c10043);
fa10044 : full_adder port map(p(447),p(478),p(509),s10044,c10044);
fa10045 : full_adder port map(p(479),p(510),p(541),s10045,c10045);
fa10046 : full_adder port map(p(511),p(542),p(573),s10046,c10046);
fa10047 : full_adder port map(p(543),p(574),p(605),s10047,c10047);
fa10048 : full_adder port map(p(575),p(606),p(637),s10048,c10048);
fa10049 : full_adder port map(p(607),p(638),p(669),s10049,c10049);
fa10050 : full_adder port map(p(639),p(670),p(701),s10050,c10050);
fa10051 : full_adder port map(p(671),p(702),p(733),s10051,c10051);
fa10052 : full_adder port map(p(703),p(734),p(765),s10052,c10052);
fa10053 : full_adder port map(p(735),p(766),p(797),s10053,c10053);
fa10054 : full_adder port map(p(767),p(798),p(829),s10054,c10054);
fa10055 : full_adder port map(p(799),p(830),p(861),s10055,c10055);
fa10056 : full_adder port map(p(831),p(862),p(893),s10056,c10056);
fa10057 : full_adder port map(p(863),p(894),p(925),s10057,c10057);
fa10058 : full_adder port map(p(895),p(926),p(957),s10058,c10058);
fa10059 : full_adder port map(p(927),p(958),p(989),s10059,c10059);
fa10060 : full_adder port map(p(959),p(990),p(1021),s10060,c10060);

--STAGE 1 GROUP 01
fa10105 : full_adder port map(p(98),p(129),p(160),s10105,c10105);
fa10106 : full_adder port map(p(99),p(130),p(161),s10106,c10106);
fa10107 : full_adder port map(p(100),p(131),p(162),s10107,c10107);
fa10108 : full_adder port map(p(101),p(132),p(163),s10108,c10108);
fa10109 : full_adder port map(p(102),p(133),p(164),s10109,c10109);
fa10110 : full_adder port map(p(103),p(134),p(165),s10110,c10110);
fa10111 : full_adder port map(p(104),p(135),p(166),s10111,c10111);
fa10112 : full_adder port map(p(105),p(136),p(167),s10112,c10112);
fa10113 : full_adder port map(p(106),p(137),p(168),s10113,c10113);
fa10114 : full_adder port map(p(107),p(138),p(169),s10114,c10114);
fa10115 : full_adder port map(p(108),p(139),p(170),s10115,c10115);
fa10116 : full_adder port map(p(109),p(140),p(171),s10116,c10116);
fa10117 : full_adder port map(p(110),p(141),p(172),s10117,c10117);
fa10118 : full_adder port map(p(111),p(142),p(173),s10118,c10118);
fa10119 : full_adder port map(p(112),p(143),p(174),s10119,c10119);
fa10120 : full_adder port map(p(113),p(144),p(175),s10120,c10120);
fa10121 : full_adder port map(p(114),p(145),p(176),s10121,c10121);
fa10122 : full_adder port map(p(115),p(146),p(177),s10122,c10122);
fa10123 : full_adder port map(p(116),p(147),p(178),s10123,c10123);
fa10124 : full_adder port map(p(117),p(148),p(179),s10124,c10124);
fa10125 : full_adder port map(p(118),p(149),p(180),s10125,c10125);
fa10126 : full_adder port map(p(119),p(150),p(181),s10126,c10126);
fa10127 : full_adder port map(p(120),p(151),p(182),s10127,c10127);
fa10128 : full_adder port map(p(121),p(152),p(183),s10128,c10128);
fa10129 : full_adder port map(p(122),p(153),p(184),s10129,c10129);
fa10130 : full_adder port map(p(123),p(154),p(185),s10130,c10130);
fa10131 : full_adder port map(p(124),p(155),p(186),s10131,c10131);
fa10132 : full_adder port map(p(156),p(187),p(218),s10132,c10132);
fa10133 : full_adder port map(p(188),p(219),p(250),s10133,c10133);
fa10134 : full_adder port map(p(220),p(251),p(282),s10134,c10134);
fa10135 : full_adder port map(p(252),p(283),p(314),s10135,c10135);
fa10136 : full_adder port map(p(284),p(315),p(346),s10136,c10136);
fa10137 : full_adder port map(p(316),p(347),p(378),s10137,c10137);
fa10138 : full_adder port map(p(348),p(379),p(410),s10138,c10138);
fa10139 : full_adder port map(p(380),p(411),p(442),s10139,c10139);
fa10140 : full_adder port map(p(412),p(443),p(474),s10140,c10140);
fa10141 : full_adder port map(p(444),p(475),p(506),s10141,c10141);
fa10142 : full_adder port map(p(476),p(507),p(538),s10142,c10142);
fa10143 : full_adder port map(p(508),p(539),p(570),s10143,c10143);
fa10144 : full_adder port map(p(540),p(571),p(602),s10144,c10144);
fa10145 : full_adder port map(p(572),p(603),p(634),s10145,c10145);
fa10146 : full_adder port map(p(604),p(635),p(666),s10146,c10146);
fa10147 : full_adder port map(p(636),p(667),p(698),s10147,c10147);
fa10148 : full_adder port map(p(668),p(699),p(730),s10148,c10148);
fa10149 : full_adder port map(p(700),p(731),p(762),s10149,c10149);
fa10150 : full_adder port map(p(732),p(763),p(794),s10150,c10150);
fa10151 : full_adder port map(p(764),p(795),p(826),s10151,c10151);
fa10152 : full_adder port map(p(796),p(827),p(858),s10152,c10152);
fa10153 : full_adder port map(p(828),p(859),p(890),s10153,c10153);
fa10154 : full_adder port map(p(860),p(891),p(922),s10154,c10154);
fa10155 : full_adder port map(p(892),p(923),p(954),s10155,c10155);
fa10156 : full_adder port map(p(924),p(955),p(986),s10156,c10156);
fa10157 : full_adder port map(p(956),p(987),p(1018),s10157,c10157);

--STAGE 1 GROUP 02
fa10208 : full_adder port map(p(194),p(225),p(256),s10208,c10208);
fa10209 : full_adder port map(p(195),p(226),p(257),s10209,c10209);
fa10210 : full_adder port map(p(196),p(227),p(258),s10210,c10210);
fa10211 : full_adder port map(p(197),p(228),p(259),s10211,c10211);
fa10212 : full_adder port map(p(198),p(229),p(260),s10212,c10212);
fa10213 : full_adder port map(p(199),p(230),p(261),s10213,c10213);
fa10214 : full_adder port map(p(200),p(231),p(262),s10214,c10214);
fa10215 : full_adder port map(p(201),p(232),p(263),s10215,c10215);
fa10216 : full_adder port map(p(202),p(233),p(264),s10216,c10216);
fa10217 : full_adder port map(p(203),p(234),p(265),s10217,c10217);
fa10218 : full_adder port map(p(204),p(235),p(266),s10218,c10218);
fa10219 : full_adder port map(p(205),p(236),p(267),s10219,c10219);
fa10220 : full_adder port map(p(206),p(237),p(268),s10220,c10220);
fa10221 : full_adder port map(p(207),p(238),p(269),s10221,c10221);
fa10222 : full_adder port map(p(208),p(239),p(270),s10222,c10222);
fa10223 : full_adder port map(p(209),p(240),p(271),s10223,c10223);
fa10224 : full_adder port map(p(210),p(241),p(272),s10224,c10224);
fa10225 : full_adder port map(p(211),p(242),p(273),s10225,c10225);
fa10226 : full_adder port map(p(212),p(243),p(274),s10226,c10226);
fa10227 : full_adder port map(p(213),p(244),p(275),s10227,c10227);
fa10228 : full_adder port map(p(214),p(245),p(276),s10228,c10228);
fa10229 : full_adder port map(p(215),p(246),p(277),s10229,c10229);
fa10230 : full_adder port map(p(216),p(247),p(278),s10230,c10230);
fa10231 : full_adder port map(p(217),p(248),p(279),s10231,c10231);
fa10232 : full_adder port map(p(249),p(280),p(311),s10232,c10232);
fa10233 : full_adder port map(p(281),p(312),p(343),s10233,c10233);
fa10234 : full_adder port map(p(313),p(344),p(375),s10234,c10234);
fa10235 : full_adder port map(p(345),p(376),p(407),s10235,c10235);
fa10236 : full_adder port map(p(377),p(408),p(439),s10236,c10236);
fa10237 : full_adder port map(p(409),p(440),p(471),s10237,c10237);
fa10238 : full_adder port map(p(441),p(472),p(503),s10238,c10238);
fa10239 : full_adder port map(p(473),p(504),p(535),s10239,c10239);
fa10240 : full_adder port map(p(505),p(536),p(567),s10240,c10240);
fa10241 : full_adder port map(p(537),p(568),p(599),s10241,c10241);
fa10242 : full_adder port map(p(569),p(600),p(631),s10242,c10242);
fa10243 : full_adder port map(p(601),p(632),p(663),s10243,c10243);
fa10244 : full_adder port map(p(633),p(664),p(695),s10244,c10244);
fa10245 : full_adder port map(p(665),p(696),p(727),s10245,c10245);
fa10246 : full_adder port map(p(697),p(728),p(759),s10246,c10246);
fa10247 : full_adder port map(p(729),p(760),p(791),s10247,c10247);
fa10248 : full_adder port map(p(761),p(792),p(823),s10248,c10248);
fa10249 : full_adder port map(p(793),p(824),p(855),s10249,c10249);
fa10250 : full_adder port map(p(825),p(856),p(887),s10250,c10250);
fa10251 : full_adder port map(p(857),p(888),p(919),s10251,c10251);
fa10252 : full_adder port map(p(889),p(920),p(951),s10252,c10252);
fa10253 : full_adder port map(p(921),p(952),p(983),s10253,c10253);
fa10254 : full_adder port map(p(953),p(984),p(1015),s10254,c10254);

--STAGE 1 GROUP 03
fa10311 : full_adder port map(p(290),p(321),p(352),s10311,c10311);
fa10312 : full_adder port map(p(291),p(322),p(353),s10312,c10312);
fa10313 : full_adder port map(p(292),p(323),p(354),s10313,c10313);
fa10314 : full_adder port map(p(293),p(324),p(355),s10314,c10314);
fa10315 : full_adder port map(p(294),p(325),p(356),s10315,c10315);
fa10316 : full_adder port map(p(295),p(326),p(357),s10316,c10316);
fa10317 : full_adder port map(p(296),p(327),p(358),s10317,c10317);
fa10318 : full_adder port map(p(297),p(328),p(359),s10318,c10318);
fa10319 : full_adder port map(p(298),p(329),p(360),s10319,c10319);
fa10320 : full_adder port map(p(299),p(330),p(361),s10320,c10320);
fa10321 : full_adder port map(p(300),p(331),p(362),s10321,c10321);
fa10322 : full_adder port map(p(301),p(332),p(363),s10322,c10322);
fa10323 : full_adder port map(p(302),p(333),p(364),s10323,c10323);
fa10324 : full_adder port map(p(303),p(334),p(365),s10324,c10324);
fa10325 : full_adder port map(p(304),p(335),p(366),s10325,c10325);
fa10326 : full_adder port map(p(305),p(336),p(367),s10326,c10326);
fa10327 : full_adder port map(p(306),p(337),p(368),s10327,c10327);
fa10328 : full_adder port map(p(307),p(338),p(369),s10328,c10328);
fa10329 : full_adder port map(p(308),p(339),p(370),s10329,c10329);
fa10330 : full_adder port map(p(309),p(340),p(371),s10330,c10330);
fa10331 : full_adder port map(p(310),p(341),p(372),s10331,c10331);
fa10332 : full_adder port map(p(342),p(373),p(404),s10332,c10332);
fa10333 : full_adder port map(p(374),p(405),p(436),s10333,c10333);
fa10334 : full_adder port map(p(406),p(437),p(468),s10334,c10334);
fa10335 : full_adder port map(p(438),p(469),p(500),s10335,c10335);
fa10336 : full_adder port map(p(470),p(501),p(532),s10336,c10336);
fa10337 : full_adder port map(p(502),p(533),p(564),s10337,c10337);
fa10338 : full_adder port map(p(534),p(565),p(596),s10338,c10338);
fa10339 : full_adder port map(p(566),p(597),p(628),s10339,c10339);
fa10340 : full_adder port map(p(598),p(629),p(660),s10340,c10340);
fa10341 : full_adder port map(p(630),p(661),p(692),s10341,c10341);
fa10342 : full_adder port map(p(662),p(693),p(724),s10342,c10342);
fa10343 : full_adder port map(p(694),p(725),p(756),s10343,c10343);
fa10344 : full_adder port map(p(726),p(757),p(788),s10344,c10344);
fa10345 : full_adder port map(p(758),p(789),p(820),s10345,c10345);
fa10346 : full_adder port map(p(790),p(821),p(852),s10346,c10346);
fa10347 : full_adder port map(p(822),p(853),p(884),s10347,c10347);
fa10348 : full_adder port map(p(854),p(885),p(916),s10348,c10348);
fa10349 : full_adder port map(p(886),p(917),p(948),s10349,c10349);
fa10350 : full_adder port map(p(918),p(949),p(980),s10350,c10350);
fa10351 : full_adder port map(p(950),p(981),p(1012),s10351,c10351);

--STAGE 1 GROUP 04
fa10414 : full_adder port map(p(386),p(417),p(448),s10414,c10414);
fa10415 : full_adder port map(p(387),p(418),p(449),s10415,c10415);
fa10416 : full_adder port map(p(388),p(419),p(450),s10416,c10416);
fa10417 : full_adder port map(p(389),p(420),p(451),s10417,c10417);
fa10418 : full_adder port map(p(390),p(421),p(452),s10418,c10418);
fa10419 : full_adder port map(p(391),p(422),p(453),s10419,c10419);
fa10420 : full_adder port map(p(392),p(423),p(454),s10420,c10420);
fa10421 : full_adder port map(p(393),p(424),p(455),s10421,c10421);
fa10422 : full_adder port map(p(394),p(425),p(456),s10422,c10422);
fa10423 : full_adder port map(p(395),p(426),p(457),s10423,c10423);
fa10424 : full_adder port map(p(396),p(427),p(458),s10424,c10424);
fa10425 : full_adder port map(p(397),p(428),p(459),s10425,c10425);
fa10426 : full_adder port map(p(398),p(429),p(460),s10426,c10426);
fa10427 : full_adder port map(p(399),p(430),p(461),s10427,c10427);
fa10428 : full_adder port map(p(400),p(431),p(462),s10428,c10428);
fa10429 : full_adder port map(p(401),p(432),p(463),s10429,c10429);
fa10430 : full_adder port map(p(402),p(433),p(464),s10430,c10430);
fa10431 : full_adder port map(p(403),p(434),p(465),s10431,c10431);
fa10432 : full_adder port map(p(435),p(466),p(497),s10432,c10432);
fa10433 : full_adder port map(p(467),p(498),p(529),s10433,c10433);
fa10434 : full_adder port map(p(499),p(530),p(561),s10434,c10434);
fa10435 : full_adder port map(p(531),p(562),p(593),s10435,c10435);
fa10436 : full_adder port map(p(563),p(594),p(625),s10436,c10436);
fa10437 : full_adder port map(p(595),p(626),p(657),s10437,c10437);
fa10438 : full_adder port map(p(627),p(658),p(689),s10438,c10438);
fa10439 : full_adder port map(p(659),p(690),p(721),s10439,c10439);
fa10440 : full_adder port map(p(691),p(722),p(753),s10440,c10440);
fa10441 : full_adder port map(p(723),p(754),p(785),s10441,c10441);
fa10442 : full_adder port map(p(755),p(786),p(817),s10442,c10442);
fa10443 : full_adder port map(p(787),p(818),p(849),s10443,c10443);
fa10444 : full_adder port map(p(819),p(850),p(881),s10444,c10444);
fa10445 : full_adder port map(p(851),p(882),p(913),s10445,c10445);
fa10446 : full_adder port map(p(883),p(914),p(945),s10446,c10446);
fa10447 : full_adder port map(p(915),p(946),p(977),s10447,c10447);
fa10448 : full_adder port map(p(947),p(978),p(1009),s10448,c10448);

--STAGE 1 GROUP 05
fa10517 : full_adder port map(p(482),p(513),p(544),s10517,c10517);
fa10518 : full_adder port map(p(483),p(514),p(545),s10518,c10518);
fa10519 : full_adder port map(p(484),p(515),p(546),s10519,c10519);
fa10520 : full_adder port map(p(485),p(516),p(547),s10520,c10520);
fa10521 : full_adder port map(p(486),p(517),p(548),s10521,c10521);
fa10522 : full_adder port map(p(487),p(518),p(549),s10522,c10522);
fa10523 : full_adder port map(p(488),p(519),p(550),s10523,c10523);
fa10524 : full_adder port map(p(489),p(520),p(551),s10524,c10524);
fa10525 : full_adder port map(p(490),p(521),p(552),s10525,c10525);
fa10526 : full_adder port map(p(491),p(522),p(553),s10526,c10526);
fa10527 : full_adder port map(p(492),p(523),p(554),s10527,c10527);
fa10528 : full_adder port map(p(493),p(524),p(555),s10528,c10528);
fa10529 : full_adder port map(p(494),p(525),p(556),s10529,c10529);
fa10530 : full_adder port map(p(495),p(526),p(557),s10530,c10530);
fa10531 : full_adder port map(p(496),p(527),p(558),s10531,c10531);
fa10532 : full_adder port map(p(528),p(559),p(590),s10532,c10532);
fa10533 : full_adder port map(p(560),p(591),p(622),s10533,c10533);
fa10534 : full_adder port map(p(592),p(623),p(654),s10534,c10534);
fa10535 : full_adder port map(p(624),p(655),p(686),s10535,c10535);
fa10536 : full_adder port map(p(656),p(687),p(718),s10536,c10536);
fa10537 : full_adder port map(p(688),p(719),p(750),s10537,c10537);
fa10538 : full_adder port map(p(720),p(751),p(782),s10538,c10538);
fa10539 : full_adder port map(p(752),p(783),p(814),s10539,c10539);
fa10540 : full_adder port map(p(784),p(815),p(846),s10540,c10540);
fa10541 : full_adder port map(p(816),p(847),p(878),s10541,c10541);
fa10542 : full_adder port map(p(848),p(879),p(910),s10542,c10542);
fa10543 : full_adder port map(p(880),p(911),p(942),s10543,c10543);
fa10544 : full_adder port map(p(912),p(943),p(974),s10544,c10544);
fa10545 : full_adder port map(p(944),p(975),p(1006),s10545,c10545);

--STAGE 1 GROUP 06
fa10620 : full_adder port map(p(578),p(609),p(640),s10620,c10620);
fa10621 : full_adder port map(p(579),p(610),p(641),s10621,c10621);
fa10622 : full_adder port map(p(580),p(611),p(642),s10622,c10622);
fa10623 : full_adder port map(p(581),p(612),p(643),s10623,c10623);
fa10624 : full_adder port map(p(582),p(613),p(644),s10624,c10624);
fa10625 : full_adder port map(p(583),p(614),p(645),s10625,c10625);
fa10626 : full_adder port map(p(584),p(615),p(646),s10626,c10626);
fa10627 : full_adder port map(p(585),p(616),p(647),s10627,c10627);
fa10628 : full_adder port map(p(586),p(617),p(648),s10628,c10628);
fa10629 : full_adder port map(p(587),p(618),p(649),s10629,c10629);
fa10630 : full_adder port map(p(588),p(619),p(650),s10630,c10630);
fa10631 : full_adder port map(p(589),p(620),p(651),s10631,c10631);
fa10632 : full_adder port map(p(621),p(652),p(683),s10632,c10632);
fa10633 : full_adder port map(p(653),p(684),p(715),s10633,c10633);
fa10634 : full_adder port map(p(685),p(716),p(747),s10634,c10634);
fa10635 : full_adder port map(p(717),p(748),p(779),s10635,c10635);
fa10636 : full_adder port map(p(749),p(780),p(811),s10636,c10636);
fa10637 : full_adder port map(p(781),p(812),p(843),s10637,c10637);
fa10638 : full_adder port map(p(813),p(844),p(875),s10638,c10638);
fa10639 : full_adder port map(p(845),p(876),p(907),s10639,c10639);
fa10640 : full_adder port map(p(877),p(908),p(939),s10640,c10640);
fa10641 : full_adder port map(p(909),p(940),p(971),s10641,c10641);
fa10642 : full_adder port map(p(941),p(972),p(1003),s10642,c10642);

--STAGE 1 GROUP 07
fa10723 : full_adder port map(p(674),p(705),p(736),s10723,c10723);
fa10724 : full_adder port map(p(675),p(706),p(737),s10724,c10724);
fa10725 : full_adder port map(p(676),p(707),p(738),s10725,c10725);
fa10726 : full_adder port map(p(677),p(708),p(739),s10726,c10726);
fa10727 : full_adder port map(p(678),p(709),p(740),s10727,c10727);
fa10728 : full_adder port map(p(679),p(710),p(741),s10728,c10728);
fa10729 : full_adder port map(p(680),p(711),p(742),s10729,c10729);
fa10730 : full_adder port map(p(681),p(712),p(743),s10730,c10730);
fa10731 : full_adder port map(p(682),p(713),p(744),s10731,c10731);
fa10732 : full_adder port map(p(714),p(745),p(776),s10732,c10732);
fa10733 : full_adder port map(p(746),p(777),p(808),s10733,c10733);
fa10734 : full_adder port map(p(778),p(809),p(840),s10734,c10734);
fa10735 : full_adder port map(p(810),p(841),p(872),s10735,c10735);
fa10736 : full_adder port map(p(842),p(873),p(904),s10736,c10736);
fa10737 : full_adder port map(p(874),p(905),p(936),s10737,c10737);
fa10738 : full_adder port map(p(906),p(937),p(968),s10738,c10738);
fa10739 : full_adder port map(p(938),p(969),p(1000),s10739,c10739);

--STAGE 1 GROUP 08
fa10826 : full_adder port map(p(770),p(801),p(832),s10826,c10826);
fa10827 : full_adder port map(p(771),p(802),p(833),s10827,c10827);
fa10828 : full_adder port map(p(772),p(803),p(834),s10828,c10828);
fa10829 : full_adder port map(p(773),p(804),p(835),s10829,c10829);
fa10830 : full_adder port map(p(774),p(805),p(836),s10830,c10830);
fa10831 : full_adder port map(p(775),p(806),p(837),s10831,c10831);
fa10832 : full_adder port map(p(807),p(838),p(869),s10832,c10832);
fa10833 : full_adder port map(p(839),p(870),p(901),s10833,c10833);
fa10834 : full_adder port map(p(871),p(902),p(933),s10834,c10834);
fa10835 : full_adder port map(p(903),p(934),p(965),s10835,c10835);
fa10836 : full_adder port map(p(935),p(966),p(997),s10836,c10836);

--STAGE 1 GROUP 09
fa10929 : full_adder port map(p(866),p(897),p(928),s10929,c10929);
fa10930 : full_adder port map(p(867),p(898),p(929),s10930,c10930);
fa10931 : full_adder port map(p(868),p(899),p(930),s10931,c10931);
fa10932 : full_adder port map(p(900),p(931),p(962),s10932,c10932);
fa10933 : full_adder port map(p(932),p(963),p(994),s10933,c10933);

-----------------------------------------------------------------

--STAGE 2 -  FULL ADDERS:214 | HALF ADDERS:0
--GROUP 00
fa20003 : full_adder port map(s10003,c10002,p(96),s20003,c20003);
fa20004 : full_adder port map(s10004,c10003,p(97),s20004,c20004);
fa20005 : full_adder port map(s10005,c10004,s10105,s20005,c20005);
fa20006 : full_adder port map(s10006,c10005,s10106,s20006,c20006);
fa20007 : full_adder port map(s10007,c10006,s10107,s20007,c20007);
fa20008 : full_adder port map(s10008,c10007,s10108,s20008,c20008);
fa20009 : full_adder port map(s10009,c10008,s10109,s20009,c20009);
fa20010 : full_adder port map(s10010,c10009,s10110,s20010,c20010);
fa20011 : full_adder port map(s10011,c10010,s10111,s20011,c20011);
fa20012 : full_adder port map(s10012,c10011,s10112,s20012,c20012);
fa20013 : full_adder port map(s10013,c10012,s10113,s20013,c20013);
fa20014 : full_adder port map(s10014,c10013,s10114,s20014,c20014);
fa20015 : full_adder port map(s10015,c10014,s10115,s20015,c20015);
fa20016 : full_adder port map(s10016,c10015,s10116,s20016,c20016);
fa20017 : full_adder port map(s10017,c10016,s10117,s20017,c20017);
fa20018 : full_adder port map(s10018,c10017,s10118,s20018,c20018);
fa20019 : full_adder port map(s10019,c10018,s10119,s20019,c20019);
fa20020 : full_adder port map(s10020,c10019,s10120,s20020,c20020);
fa20021 : full_adder port map(s10021,c10020,s10121,s20021,c20021);
fa20022 : full_adder port map(s10022,c10021,s10122,s20022,c20022);
fa20023 : full_adder port map(s10023,c10022,s10123,s20023,c20023);
fa20024 : full_adder port map(s10024,c10023,s10124,s20024,c20024);
fa20025 : full_adder port map(s10025,c10024,s10125,s20025,c20025);
fa20026 : full_adder port map(s10026,c10025,s10126,s20026,c20026);
fa20027 : full_adder port map(s10027,c10026,s10127,s20027,c20027);
fa20028 : full_adder port map(s10028,c10027,s10128,s20028,c20028);
fa20029 : full_adder port map(s10029,c10028,s10129,s20029,c20029);
fa20030 : full_adder port map(s10030,c10029,s10130,s20030,c20030);
fa20031 : full_adder port map(s10031,c10030,s10131,s20031,c20031);
fa20032 : full_adder port map(s10032,c10031,s10132,s20032,c20032);
fa20033 : full_adder port map(s10033,c10032,s10133,s20033,c20033);
fa20034 : full_adder port map(s10034,c10033,s10134,s20034,c20034);
fa20035 : full_adder port map(s10035,c10034,s10135,s20035,c20035);
fa20036 : full_adder port map(s10036,c10035,s10136,s20036,c20036);
fa20037 : full_adder port map(s10037,c10036,s10137,s20037,c20037);
fa20038 : full_adder port map(s10038,c10037,s10138,s20038,c20038);
fa20039 : full_adder port map(s10039,c10038,s10139,s20039,c20039);
fa20040 : full_adder port map(s10040,c10039,s10140,s20040,c20040);
fa20041 : full_adder port map(s10041,c10040,s10141,s20041,c20041);
fa20042 : full_adder port map(s10042,c10041,s10142,s20042,c20042);
fa20043 : full_adder port map(s10043,c10042,s10143,s20043,c20043);
fa20044 : full_adder port map(s10044,c10043,s10144,s20044,c20044);
fa20045 : full_adder port map(s10045,c10044,s10145,s20045,c20045);
fa20046 : full_adder port map(s10046,c10045,s10146,s20046,c20046);
fa20047 : full_adder port map(s10047,c10046,s10147,s20047,c20047);
fa20048 : full_adder port map(s10048,c10047,s10148,s20048,c20048);
fa20049 : full_adder port map(s10049,c10048,s10149,s20049,c20049);
fa20050 : full_adder port map(s10050,c10049,s10150,s20050,c20050);
fa20051 : full_adder port map(s10051,c10050,s10151,s20051,c20051);
fa20052 : full_adder port map(s10052,c10051,s10152,s20052,c20052);
fa20053 : full_adder port map(s10053,c10052,s10153,s20053,c20053);
fa20054 : full_adder port map(s10054,c10053,s10154,s20054,c20054);
fa20055 : full_adder port map(s10055,c10054,s10155,s20055,c20055);
fa20056 : full_adder port map(s10056,c10055,s10156,s20056,c20056);
fa20057 : full_adder port map(s10057,c10056,s10157,s20057,c20057);
fa20058 : full_adder port map(s10058,c10057,p(988),s20058,c20058);
fa20059 : full_adder port map(s10059,c10058,p(1020),s20059,c20059);
fa20061 : full_adder port map(p(991),p(1022),c10060,s20061,c20061);

--STAGE 2 GROUP 01
fa20107 : full_adder port map(c10106,p(193),p(224),s20107,c20107);
fa20109 : full_adder port map(c10108,s10209,c10208,s20109,c20109);
fa20110 : full_adder port map(c10109,s10210,c10209,s20110,c20110);
fa20111 : full_adder port map(c10110,s10211,c10210,s20111,c20111);
fa20112 : full_adder port map(c10111,s10212,c10211,s20112,c20112);
fa20113 : full_adder port map(c10112,s10213,c10212,s20113,c20113);
fa20114 : full_adder port map(c10113,s10214,c10213,s20114,c20114);
fa20115 : full_adder port map(c10114,s10215,c10214,s20115,c20115);
fa20116 : full_adder port map(c10115,s10216,c10215,s20116,c20116);
fa20117 : full_adder port map(c10116,s10217,c10216,s20117,c20117);
fa20118 : full_adder port map(c10117,s10218,c10217,s20118,c20118);
fa20119 : full_adder port map(c10118,s10219,c10218,s20119,c20119);
fa20120 : full_adder port map(c10119,s10220,c10219,s20120,c20120);
fa20121 : full_adder port map(c10120,s10221,c10220,s20121,c20121);
fa20122 : full_adder port map(c10121,s10222,c10221,s20122,c20122);
fa20123 : full_adder port map(c10122,s10223,c10222,s20123,c20123);
fa20124 : full_adder port map(c10123,s10224,c10223,s20124,c20124);
fa20125 : full_adder port map(c10124,s10225,c10224,s20125,c20125);
fa20126 : full_adder port map(c10125,s10226,c10225,s20126,c20126);
fa20127 : full_adder port map(c10126,s10227,c10226,s20127,c20127);
fa20128 : full_adder port map(c10127,s10228,c10227,s20128,c20128);
fa20129 : full_adder port map(c10128,s10229,c10228,s20129,c20129);
fa20130 : full_adder port map(c10129,s10230,c10229,s20130,c20130);
fa20131 : full_adder port map(c10130,s10231,c10230,s20131,c20131);
fa20132 : full_adder port map(c10131,s10232,c10231,s20132,c20132);
fa20133 : full_adder port map(c10132,s10233,c10232,s20133,c20133);
fa20134 : full_adder port map(c10133,s10234,c10233,s20134,c20134);
fa20135 : full_adder port map(c10134,s10235,c10234,s20135,c20135);
fa20136 : full_adder port map(c10135,s10236,c10235,s20136,c20136);
fa20137 : full_adder port map(c10136,s10237,c10236,s20137,c20137);
fa20138 : full_adder port map(c10137,s10238,c10237,s20138,c20138);
fa20139 : full_adder port map(c10138,s10239,c10238,s20139,c20139);
fa20140 : full_adder port map(c10139,s10240,c10239,s20140,c20140);
fa20141 : full_adder port map(c10140,s10241,c10240,s20141,c20141);
fa20142 : full_adder port map(c10141,s10242,c10241,s20142,c20142);
fa20143 : full_adder port map(c10142,s10243,c10242,s20143,c20143);
fa20144 : full_adder port map(c10143,s10244,c10243,s20144,c20144);
fa20145 : full_adder port map(c10144,s10245,c10244,s20145,c20145);
fa20146 : full_adder port map(c10145,s10246,c10245,s20146,c20146);
fa20147 : full_adder port map(c10146,s10247,c10246,s20147,c20147);
fa20148 : full_adder port map(c10147,s10248,c10247,s20148,c20148);
fa20149 : full_adder port map(c10148,s10249,c10248,s20149,c20149);
fa20150 : full_adder port map(c10149,s10250,c10249,s20150,c20150);
fa20151 : full_adder port map(c10150,s10251,c10250,s20151,c20151);
fa20152 : full_adder port map(c10151,s10252,c10251,s20152,c20152);
fa20153 : full_adder port map(c10152,s10253,c10252,s20153,c20153);
fa20154 : full_adder port map(c10153,s10254,c10253,s20154,c20154);
fa20155 : full_adder port map(c10154,p(985),p(1016),s20155,c20155);

--STAGE 2 GROUP 02
fa20212 : full_adder port map(s10312,c10311,p(384),s20212,c20212);
fa20213 : full_adder port map(s10313,c10312,p(385),s20213,c20213);
fa20214 : full_adder port map(s10314,c10313,s10414,s20214,c20214);
fa20215 : full_adder port map(s10315,c10314,s10415,s20215,c20215);
fa20216 : full_adder port map(s10316,c10315,s10416,s20216,c20216);
fa20217 : full_adder port map(s10317,c10316,s10417,s20217,c20217);
fa20218 : full_adder port map(s10318,c10317,s10418,s20218,c20218);
fa20219 : full_adder port map(s10319,c10318,s10419,s20219,c20219);
fa20220 : full_adder port map(s10320,c10319,s10420,s20220,c20220);
fa20221 : full_adder port map(s10321,c10320,s10421,s20221,c20221);
fa20222 : full_adder port map(s10322,c10321,s10422,s20222,c20222);
fa20223 : full_adder port map(s10323,c10322,s10423,s20223,c20223);
fa20224 : full_adder port map(s10324,c10323,s10424,s20224,c20224);
fa20225 : full_adder port map(s10325,c10324,s10425,s20225,c20225);
fa20226 : full_adder port map(s10326,c10325,s10426,s20226,c20226);
fa20227 : full_adder port map(s10327,c10326,s10427,s20227,c20227);
fa20228 : full_adder port map(s10328,c10327,s10428,s20228,c20228);
fa20229 : full_adder port map(s10329,c10328,s10429,s20229,c20229);
fa20230 : full_adder port map(s10330,c10329,s10430,s20230,c20230);
fa20231 : full_adder port map(s10331,c10330,s10431,s20231,c20231);
fa20232 : full_adder port map(s10332,c10331,s10432,s20232,c20232);
fa20233 : full_adder port map(s10333,c10332,s10433,s20233,c20233);
fa20234 : full_adder port map(s10334,c10333,s10434,s20234,c20234);
fa20235 : full_adder port map(s10335,c10334,s10435,s20235,c20235);
fa20236 : full_adder port map(s10336,c10335,s10436,s20236,c20236);
fa20237 : full_adder port map(s10337,c10336,s10437,s20237,c20237);
fa20238 : full_adder port map(s10338,c10337,s10438,s20238,c20238);
fa20239 : full_adder port map(s10339,c10338,s10439,s20239,c20239);
fa20240 : full_adder port map(s10340,c10339,s10440,s20240,c20240);
fa20241 : full_adder port map(s10341,c10340,s10441,s20241,c20241);
fa20242 : full_adder port map(s10342,c10341,s10442,s20242,c20242);
fa20243 : full_adder port map(s10343,c10342,s10443,s20243,c20243);
fa20244 : full_adder port map(s10344,c10343,s10444,s20244,c20244);
fa20245 : full_adder port map(s10345,c10344,s10445,s20245,c20245);
fa20246 : full_adder port map(s10346,c10345,s10446,s20246,c20246);
fa20247 : full_adder port map(s10347,c10346,s10447,s20247,c20247);
fa20248 : full_adder port map(s10348,c10347,s10448,s20248,c20248);
fa20249 : full_adder port map(s10349,c10348,p(979),s20249,c20249);
fa20250 : full_adder port map(s10350,c10349,p(1011),s20250,c20250);
fa20252 : full_adder port map(p(982),p(1013),c10351,s20252,c20252);

--STAGE 2 GROUP 03
fa20316 : full_adder port map(c10415,p(481),p(512),s20316,c20316);
fa20318 : full_adder port map(c10417,s10518,c10517,s20318,c20318);
fa20319 : full_adder port map(c10418,s10519,c10518,s20319,c20319);
fa20320 : full_adder port map(c10419,s10520,c10519,s20320,c20320);
fa20321 : full_adder port map(c10420,s10521,c10520,s20321,c20321);
fa20322 : full_adder port map(c10421,s10522,c10521,s20322,c20322);
fa20323 : full_adder port map(c10422,s10523,c10522,s20323,c20323);
fa20324 : full_adder port map(c10423,s10524,c10523,s20324,c20324);
fa20325 : full_adder port map(c10424,s10525,c10524,s20325,c20325);
fa20326 : full_adder port map(c10425,s10526,c10525,s20326,c20326);
fa20327 : full_adder port map(c10426,s10527,c10526,s20327,c20327);
fa20328 : full_adder port map(c10427,s10528,c10527,s20328,c20328);
fa20329 : full_adder port map(c10428,s10529,c10528,s20329,c20329);
fa20330 : full_adder port map(c10429,s10530,c10529,s20330,c20330);
fa20331 : full_adder port map(c10430,s10531,c10530,s20331,c20331);
fa20332 : full_adder port map(c10431,s10532,c10531,s20332,c20332);
fa20333 : full_adder port map(c10432,s10533,c10532,s20333,c20333);
fa20334 : full_adder port map(c10433,s10534,c10533,s20334,c20334);
fa20335 : full_adder port map(c10434,s10535,c10534,s20335,c20335);
fa20336 : full_adder port map(c10435,s10536,c10535,s20336,c20336);
fa20337 : full_adder port map(c10436,s10537,c10536,s20337,c20337);
fa20338 : full_adder port map(c10437,s10538,c10537,s20338,c20338);
fa20339 : full_adder port map(c10438,s10539,c10538,s20339,c20339);
fa20340 : full_adder port map(c10439,s10540,c10539,s20340,c20340);
fa20341 : full_adder port map(c10440,s10541,c10540,s20341,c20341);
fa20342 : full_adder port map(c10441,s10542,c10541,s20342,c20342);
fa20343 : full_adder port map(c10442,s10543,c10542,s20343,c20343);
fa20344 : full_adder port map(c10443,s10544,c10543,s20344,c20344);
fa20345 : full_adder port map(c10444,s10545,c10544,s20345,c20345);
fa20346 : full_adder port map(c10445,p(976),p(1007),s20346,c20346);

--STAGE 2 GROUP 04
fa20421 : full_adder port map(s10621,c10620,p(672),s20421,c20421);
fa20422 : full_adder port map(s10622,c10621,p(673),s20422,c20422);
fa20423 : full_adder port map(s10623,c10622,s10723,s20423,c20423);
fa20424 : full_adder port map(s10624,c10623,s10724,s20424,c20424);
fa20425 : full_adder port map(s10625,c10624,s10725,s20425,c20425);
fa20426 : full_adder port map(s10626,c10625,s10726,s20426,c20426);
fa20427 : full_adder port map(s10627,c10626,s10727,s20427,c20427);
fa20428 : full_adder port map(s10628,c10627,s10728,s20428,c20428);
fa20429 : full_adder port map(s10629,c10628,s10729,s20429,c20429);
fa20430 : full_adder port map(s10630,c10629,s10730,s20430,c20430);
fa20431 : full_adder port map(s10631,c10630,s10731,s20431,c20431);
fa20432 : full_adder port map(s10632,c10631,s10732,s20432,c20432);
fa20433 : full_adder port map(s10633,c10632,s10733,s20433,c20433);
fa20434 : full_adder port map(s10634,c10633,s10734,s20434,c20434);
fa20435 : full_adder port map(s10635,c10634,s10735,s20435,c20435);
fa20436 : full_adder port map(s10636,c10635,s10736,s20436,c20436);
fa20437 : full_adder port map(s10637,c10636,s10737,s20437,c20437);
fa20438 : full_adder port map(s10638,c10637,s10738,s20438,c20438);
fa20439 : full_adder port map(s10639,c10638,s10739,s20439,c20439);
fa20440 : full_adder port map(s10640,c10639,p(970),s20440,c20440);
fa20441 : full_adder port map(s10641,c10640,p(1002),s20441,c20441);
fa20443 : full_adder port map(p(973),p(1004),c10642,s20443,c20443);

--STAGE 2 GROUP 05
fa20525 : full_adder port map(c10724,p(769),p(800),s20525,c20525);
fa20527 : full_adder port map(c10726,s10827,c10826,s20527,c20527);
fa20528 : full_adder port map(c10727,s10828,c10827,s20528,c20528);
fa20529 : full_adder port map(c10728,s10829,c10828,s20529,c20529);
fa20530 : full_adder port map(c10729,s10830,c10829,s20530,c20530);
fa20531 : full_adder port map(c10730,s10831,c10830,s20531,c20531);
fa20532 : full_adder port map(c10731,s10832,c10831,s20532,c20532);
fa20533 : full_adder port map(c10732,s10833,c10832,s20533,c20533);
fa20534 : full_adder port map(c10733,s10834,c10833,s20534,c20534);
fa20535 : full_adder port map(c10734,s10835,c10834,s20535,c20535);
fa20536 : full_adder port map(c10735,s10836,c10835,s20536,c20536);
fa20537 : full_adder port map(c10736,p(967),p(998),s20537,c20537);

--STAGE 2 GROUP 06
fa20630 : full_adder port map(s10930,c10929,p(960),s20630,c20630);
fa20631 : full_adder port map(s10931,c10930,p(961),s20631,c20631);
fa20632 : full_adder port map(s10932,c10931,p(993),s20632,c20632);
fa20634 : full_adder port map(p(964),p(995),c10933,s20634,c20634);

-----------------------------------------------------------------

--STAGE 3 -  FULL ADDERS:142 | HALF ADDERS:19
--GROUP 00
fa30004 : full_adder port map(s20004,c20003,p(128),s30004,c30004);
ha30005 : half_adder port map(s20005,c20004,s30005,c30005);
fa30006 : full_adder port map(s20006,c20005,c10105,s30006,c30006);
fa30007 : full_adder port map(s20007,c20006,s20107,s30007,c30007);
fa30008 : full_adder port map(s20008,c20007,c10107,s30008,c30008);
fa30009 : full_adder port map(s20009,c20008,s20109,s30009,c30009);
fa30010 : full_adder port map(s20010,c20009,s20110,s30010,c30010);
fa30011 : full_adder port map(s20011,c20010,s20111,s30011,c30011);
fa30012 : full_adder port map(s20012,c20011,s20112,s30012,c30012);
fa30013 : full_adder port map(s20013,c20012,s20113,s30013,c30013);
fa30014 : full_adder port map(s20014,c20013,s20114,s30014,c30014);
fa30015 : full_adder port map(s20015,c20014,s20115,s30015,c30015);
fa30016 : full_adder port map(s20016,c20015,s20116,s30016,c30016);
fa30017 : full_adder port map(s20017,c20016,s20117,s30017,c30017);
fa30018 : full_adder port map(s20018,c20017,s20118,s30018,c30018);
fa30019 : full_adder port map(s20019,c20018,s20119,s30019,c30019);
fa30020 : full_adder port map(s20020,c20019,s20120,s30020,c30020);
fa30021 : full_adder port map(s20021,c20020,s20121,s30021,c30021);
fa30022 : full_adder port map(s20022,c20021,s20122,s30022,c30022);
fa30023 : full_adder port map(s20023,c20022,s20123,s30023,c30023);
fa30024 : full_adder port map(s20024,c20023,s20124,s30024,c30024);
fa30025 : full_adder port map(s20025,c20024,s20125,s30025,c30025);
fa30026 : full_adder port map(s20026,c20025,s20126,s30026,c30026);
fa30027 : full_adder port map(s20027,c20026,s20127,s30027,c30027);
fa30028 : full_adder port map(s20028,c20027,s20128,s30028,c30028);
fa30029 : full_adder port map(s20029,c20028,s20129,s30029,c30029);
fa30030 : full_adder port map(s20030,c20029,s20130,s30030,c30030);
fa30031 : full_adder port map(s20031,c20030,s20131,s30031,c30031);
fa30032 : full_adder port map(s20032,c20031,s20132,s30032,c30032);
fa30033 : full_adder port map(s20033,c20032,s20133,s30033,c30033);
fa30034 : full_adder port map(s20034,c20033,s20134,s30034,c30034);
fa30035 : full_adder port map(s20035,c20034,s20135,s30035,c30035);
fa30036 : full_adder port map(s20036,c20035,s20136,s30036,c30036);
fa30037 : full_adder port map(s20037,c20036,s20137,s30037,c30037);
fa30038 : full_adder port map(s20038,c20037,s20138,s30038,c30038);
fa30039 : full_adder port map(s20039,c20038,s20139,s30039,c30039);
fa30040 : full_adder port map(s20040,c20039,s20140,s30040,c30040);
fa30041 : full_adder port map(s20041,c20040,s20141,s30041,c30041);
fa30042 : full_adder port map(s20042,c20041,s20142,s30042,c30042);
fa30043 : full_adder port map(s20043,c20042,s20143,s30043,c30043);
fa30044 : full_adder port map(s20044,c20043,s20144,s30044,c30044);
fa30045 : full_adder port map(s20045,c20044,s20145,s30045,c30045);
fa30046 : full_adder port map(s20046,c20045,s20146,s30046,c30046);
fa30047 : full_adder port map(s20047,c20046,s20147,s30047,c30047);
fa30048 : full_adder port map(s20048,c20047,s20148,s30048,c30048);
fa30049 : full_adder port map(s20049,c20048,s20149,s30049,c30049);
fa30050 : full_adder port map(s20050,c20049,s20150,s30050,c30050);
fa30051 : full_adder port map(s20051,c20050,s20151,s30051,c30051);
fa30052 : full_adder port map(s20052,c20051,s20152,s30052,c30052);
fa30053 : full_adder port map(s20053,c20052,s20153,s30053,c30053);
fa30054 : full_adder port map(s20054,c20053,s20154,s30054,c30054);
fa30055 : full_adder port map(s20055,c20054,s20155,s30055,c30055);
fa30056 : full_adder port map(s20056,c20055,c10155,s30056,c30056);
fa30057 : full_adder port map(s20057,c20056,c10156,s30057,c30057);
fa30058 : full_adder port map(s20058,c20057,p(1019),s30058,c30058);
ha30059 : half_adder port map(s20059,c20058,s30059,c30059);
fa30060 : full_adder port map(s10060,c10059,c20059,s30060,c30060);

--STAGE 3 GROUP 01
ha30108 : half_adder port map(s10208,c20107,s30108,c30108);
fa30110 : full_adder port map(c20109,p(289),p(320),s30110,c30110);
ha30111 : half_adder port map(c20110,s10311,s30111,c30111);
ha30112 : half_adder port map(c20111,s20212,s30112,c30112);
fa30113 : full_adder port map(c20112,s20213,c20212,s30113,c30113);
fa30114 : full_adder port map(c20113,s20214,c20213,s30114,c30114);
fa30115 : full_adder port map(c20114,s20215,c20214,s30115,c30115);
fa30116 : full_adder port map(c20115,s20216,c20215,s30116,c30116);
fa30117 : full_adder port map(c20116,s20217,c20216,s30117,c30117);
fa30118 : full_adder port map(c20117,s20218,c20217,s30118,c30118);
fa30119 : full_adder port map(c20118,s20219,c20218,s30119,c30119);
fa30120 : full_adder port map(c20119,s20220,c20219,s30120,c30120);
fa30121 : full_adder port map(c20120,s20221,c20220,s30121,c30121);
fa30122 : full_adder port map(c20121,s20222,c20221,s30122,c30122);
fa30123 : full_adder port map(c20122,s20223,c20222,s30123,c30123);
fa30124 : full_adder port map(c20123,s20224,c20223,s30124,c30124);
fa30125 : full_adder port map(c20124,s20225,c20224,s30125,c30125);
fa30126 : full_adder port map(c20125,s20226,c20225,s30126,c30126);
fa30127 : full_adder port map(c20126,s20227,c20226,s30127,c30127);
fa30128 : full_adder port map(c20127,s20228,c20227,s30128,c30128);
fa30129 : full_adder port map(c20128,s20229,c20228,s30129,c30129);
fa30130 : full_adder port map(c20129,s20230,c20229,s30130,c30130);
fa30131 : full_adder port map(c20130,s20231,c20230,s30131,c30131);
fa30132 : full_adder port map(c20131,s20232,c20231,s30132,c30132);
fa30133 : full_adder port map(c20132,s20233,c20232,s30133,c30133);
fa30134 : full_adder port map(c20133,s20234,c20233,s30134,c30134);
fa30135 : full_adder port map(c20134,s20235,c20234,s30135,c30135);
fa30136 : full_adder port map(c20135,s20236,c20235,s30136,c30136);
fa30137 : full_adder port map(c20136,s20237,c20236,s30137,c30137);
fa30138 : full_adder port map(c20137,s20238,c20237,s30138,c30138);
fa30139 : full_adder port map(c20138,s20239,c20238,s30139,c30139);
fa30140 : full_adder port map(c20139,s20240,c20239,s30140,c30140);
fa30141 : full_adder port map(c20140,s20241,c20240,s30141,c30141);
fa30142 : full_adder port map(c20141,s20242,c20241,s30142,c30142);
fa30143 : full_adder port map(c20142,s20243,c20242,s30143,c30143);
fa30144 : full_adder port map(c20143,s20244,c20243,s30144,c30144);
fa30145 : full_adder port map(c20144,s20245,c20244,s30145,c30145);
fa30146 : full_adder port map(c20145,s20246,c20245,s30146,c30146);
fa30147 : full_adder port map(c20146,s20247,c20246,s30147,c30147);
fa30148 : full_adder port map(c20147,s20248,c20247,s30148,c30148);
fa30149 : full_adder port map(c20148,s20249,c20248,s30149,c30149);
fa30150 : full_adder port map(c20149,s20250,c20249,s30150,c30150);
fa30151 : full_adder port map(c20150,s10351,c10350,s30151,c30151);
ha30152 : half_adder port map(c20151,s20252,s30152,c30152);
fa30153 : full_adder port map(c20152,p(1014),c20252,s30153,c30153);
ha30155 : half_adder port map(c20154,c10254,s30155,c30155);
ha30156 : half_adder port map(p(1017),c20155,s30156,c30156);

--STAGE 3 GROUP 02
ha30215 : half_adder port map(c10414,p(480),s30215,c30215);
fa30217 : full_adder port map(c10416,s10517,c20316,s30217,c30217);
ha30218 : half_adder port map(s20318,p(576),s30218,c30218);
fa30219 : full_adder port map(s20319,c20318,p(577),s30219,c30219);
fa30220 : full_adder port map(s20320,c20319,s10620,s30220,c30220);
fa30221 : full_adder port map(s20321,c20320,s20421,s30221,c30221);
fa30222 : full_adder port map(s20322,c20321,s20422,s30222,c30222);
fa30223 : full_adder port map(s20323,c20322,s20423,s30223,c30223);
fa30224 : full_adder port map(s20324,c20323,s20424,s30224,c30224);
fa30225 : full_adder port map(s20325,c20324,s20425,s30225,c30225);
fa30226 : full_adder port map(s20326,c20325,s20426,s30226,c30226);
fa30227 : full_adder port map(s20327,c20326,s20427,s30227,c30227);
fa30228 : full_adder port map(s20328,c20327,s20428,s30228,c30228);
fa30229 : full_adder port map(s20329,c20328,s20429,s30229,c30229);
fa30230 : full_adder port map(s20330,c20329,s20430,s30230,c30230);
fa30231 : full_adder port map(s20331,c20330,s20431,s30231,c30231);
fa30232 : full_adder port map(s20332,c20331,s20432,s30232,c30232);
fa30233 : full_adder port map(s20333,c20332,s20433,s30233,c30233);
fa30234 : full_adder port map(s20334,c20333,s20434,s30234,c30234);
fa30235 : full_adder port map(s20335,c20334,s20435,s30235,c30235);
fa30236 : full_adder port map(s20336,c20335,s20436,s30236,c30236);
fa30237 : full_adder port map(s20337,c20336,s20437,s30237,c30237);
fa30238 : full_adder port map(s20338,c20337,s20438,s30238,c30238);
fa30239 : full_adder port map(s20339,c20338,s20439,s30239,c30239);
fa30240 : full_adder port map(s20340,c20339,s20440,s30240,c30240);
fa30241 : full_adder port map(s20341,c20340,s20441,s30241,c30241);
fa30242 : full_adder port map(s20342,c20341,s10642,s30242,c30242);
fa30243 : full_adder port map(s20343,c20342,s20443,s30243,c30243);
fa30244 : full_adder port map(s20344,c20343,p(1005),s30244,c30244);
ha30245 : half_adder port map(s20345,c20344,s30245,c30245);
fa30246 : full_adder port map(s20346,c20345,c10545,s30246,c30246);
fa30247 : full_adder port map(c10446,p(1008),c20346,s30247,c30247);
ha30249 : half_adder port map(p(1010),c10448,s30249,c30249);

--STAGE 3 GROUP 03
ha30322 : half_adder port map(c20421,p(704),s30322,c30322);
fa30324 : full_adder port map(c20423,c10723,p(768),s30324,c30324);
ha30325 : half_adder port map(c20424,s20525,s30325,c30325);
fa30326 : full_adder port map(c20425,c10725,s10826,s30326,c30326);
fa30327 : full_adder port map(c20426,s20527,p(864),s30327,c30327);
fa30328 : full_adder port map(c20427,s20528,c20527,s30328,c30328);
fa30329 : full_adder port map(c20428,s20529,c20528,s30329,c30329);
fa30330 : full_adder port map(c20429,s20530,c20529,s30330,c30330);
fa30331 : full_adder port map(c20430,s20531,c20530,s30331,c30331);
fa30332 : full_adder port map(c20431,s20532,c20531,s30332,c30332);
fa30333 : full_adder port map(c20432,s20533,c20532,s30333,c30333);
fa30334 : full_adder port map(c20433,s20534,c20533,s30334,c30334);
fa30335 : full_adder port map(c20434,s20535,c20534,s30335,c30335);
fa30336 : full_adder port map(c20435,s20536,c20535,s30336,c30336);
fa30337 : full_adder port map(c20436,s20537,c20536,s30337,c30337);
fa30338 : full_adder port map(c20437,c10737,p(999),s30338,c30338);
ha30339 : half_adder port map(c20438,c10738,s30339,c30339);
fa30340 : full_adder port map(c20439,p(1001),c10739,s30340,c30340);
ha30342 : half_adder port map(c10641,c20441,s30342,c30342);

--STAGE 3 GROUP 04
ha30428 : half_adder port map(p(865),p(896),s30428,c30428);
fa30431 : full_adder port map(s20631,c20630,p(992),s30431,c30431);
ha30432 : half_adder port map(s20632,c20631,s30432,c30432);
fa30433 : full_adder port map(s10933,c10932,c20632,s30433,c30433);
ha30435 : half_adder port map(p(996),c20634,s30435,c30435);

-----------------------------------------------------------------

--STAGE 4 -  FULL ADDERS:96 | HALF ADDERS:0
--GROUP 00
fa40006 : full_adder port map(s30006,c30005,p(192),s40006,c40006);
fa40008 : full_adder port map(s30008,c30007,s30108,s40008,c40008);
fa40009 : full_adder port map(s30009,c30008,p(288),s40009,c40009);
fa40010 : full_adder port map(s30010,c30009,s30110,s40010,c40010);
fa40011 : full_adder port map(s30011,c30010,s30111,s40011,c40011);
fa40012 : full_adder port map(s30012,c30011,s30112,s40012,c40012);
fa40013 : full_adder port map(s30013,c30012,s30113,s40013,c40013);
fa40014 : full_adder port map(s30014,c30013,s30114,s40014,c40014);
fa40015 : full_adder port map(s30015,c30014,s30115,s40015,c40015);
fa40016 : full_adder port map(s30016,c30015,s30116,s40016,c40016);
fa40017 : full_adder port map(s30017,c30016,s30117,s40017,c40017);
fa40018 : full_adder port map(s30018,c30017,s30118,s40018,c40018);
fa40019 : full_adder port map(s30019,c30018,s30119,s40019,c40019);
fa40020 : full_adder port map(s30020,c30019,s30120,s40020,c40020);
fa40021 : full_adder port map(s30021,c30020,s30121,s40021,c40021);
fa40022 : full_adder port map(s30022,c30021,s30122,s40022,c40022);
fa40023 : full_adder port map(s30023,c30022,s30123,s40023,c40023);
fa40024 : full_adder port map(s30024,c30023,s30124,s40024,c40024);
fa40025 : full_adder port map(s30025,c30024,s30125,s40025,c40025);
fa40026 : full_adder port map(s30026,c30025,s30126,s40026,c40026);
fa40027 : full_adder port map(s30027,c30026,s30127,s40027,c40027);
fa40028 : full_adder port map(s30028,c30027,s30128,s40028,c40028);
fa40029 : full_adder port map(s30029,c30028,s30129,s40029,c40029);
fa40030 : full_adder port map(s30030,c30029,s30130,s40030,c40030);
fa40031 : full_adder port map(s30031,c30030,s30131,s40031,c40031);
fa40032 : full_adder port map(s30032,c30031,s30132,s40032,c40032);
fa40033 : full_adder port map(s30033,c30032,s30133,s40033,c40033);
fa40034 : full_adder port map(s30034,c30033,s30134,s40034,c40034);
fa40035 : full_adder port map(s30035,c30034,s30135,s40035,c40035);
fa40036 : full_adder port map(s30036,c30035,s30136,s40036,c40036);
fa40037 : full_adder port map(s30037,c30036,s30137,s40037,c40037);
fa40038 : full_adder port map(s30038,c30037,s30138,s40038,c40038);
fa40039 : full_adder port map(s30039,c30038,s30139,s40039,c40039);
fa40040 : full_adder port map(s30040,c30039,s30140,s40040,c40040);
fa40041 : full_adder port map(s30041,c30040,s30141,s40041,c40041);
fa40042 : full_adder port map(s30042,c30041,s30142,s40042,c40042);
fa40043 : full_adder port map(s30043,c30042,s30143,s40043,c40043);
fa40044 : full_adder port map(s30044,c30043,s30144,s40044,c40044);
fa40045 : full_adder port map(s30045,c30044,s30145,s40045,c40045);
fa40046 : full_adder port map(s30046,c30045,s30146,s40046,c40046);
fa40047 : full_adder port map(s30047,c30046,s30147,s40047,c40047);
fa40048 : full_adder port map(s30048,c30047,s30148,s40048,c40048);
fa40049 : full_adder port map(s30049,c30048,s30149,s40049,c40049);
fa40050 : full_adder port map(s30050,c30049,s30150,s40050,c40050);
fa40051 : full_adder port map(s30051,c30050,s30151,s40051,c40051);
fa40052 : full_adder port map(s30052,c30051,s30152,s40052,c40052);
fa40053 : full_adder port map(s30053,c30052,s30153,s40053,c40053);
fa40054 : full_adder port map(s30054,c30053,c20153,s40054,c40054);
fa40055 : full_adder port map(s30055,c30054,s30155,s40055,c40055);
fa40056 : full_adder port map(s30056,c30055,s30156,s40056,c40056);
fa40057 : full_adder port map(s30057,c30056,c30156,s40057,c40057);
fa40058 : full_adder port map(s30058,c30057,c10157,s40058,c40058);

--STAGE 4 GROUP 01
fa40116 : full_adder port map(c30115,s20316,c30215,s40116,c40116);
fa40118 : full_adder port map(c30117,s30218,c30217,s40118,c40118);
fa40119 : full_adder port map(c30118,s30219,c30218,s40119,c40119);
fa40120 : full_adder port map(c30119,s30220,c30219,s40120,c40120);
fa40121 : full_adder port map(c30120,s30221,c30220,s40121,c40121);
fa40122 : full_adder port map(c30121,s30222,c30221,s40122,c40122);
fa40123 : full_adder port map(c30122,s30223,c30222,s40123,c40123);
fa40124 : full_adder port map(c30123,s30224,c30223,s40124,c40124);
fa40125 : full_adder port map(c30124,s30225,c30224,s40125,c40125);
fa40126 : full_adder port map(c30125,s30226,c30225,s40126,c40126);
fa40127 : full_adder port map(c30126,s30227,c30226,s40127,c40127);
fa40128 : full_adder port map(c30127,s30228,c30227,s40128,c40128);
fa40129 : full_adder port map(c30128,s30229,c30228,s40129,c40129);
fa40130 : full_adder port map(c30129,s30230,c30229,s40130,c40130);
fa40131 : full_adder port map(c30130,s30231,c30230,s40131,c40131);
fa40132 : full_adder port map(c30131,s30232,c30231,s40132,c40132);
fa40133 : full_adder port map(c30132,s30233,c30232,s40133,c40133);
fa40134 : full_adder port map(c30133,s30234,c30233,s40134,c40134);
fa40135 : full_adder port map(c30134,s30235,c30234,s40135,c40135);
fa40136 : full_adder port map(c30135,s30236,c30235,s40136,c40136);
fa40137 : full_adder port map(c30136,s30237,c30236,s40137,c40137);
fa40138 : full_adder port map(c30137,s30238,c30237,s40138,c40138);
fa40139 : full_adder port map(c30138,s30239,c30238,s40139,c40139);
fa40140 : full_adder port map(c30139,s30240,c30239,s40140,c40140);
fa40141 : full_adder port map(c30140,s30241,c30240,s40141,c40141);
fa40142 : full_adder port map(c30141,s30242,c30241,s40142,c40142);
fa40143 : full_adder port map(c30142,s30243,c30242,s40143,c40143);
fa40144 : full_adder port map(c30143,s30244,c30243,s40144,c40144);
fa40145 : full_adder port map(c30144,s30245,c30244,s40145,c40145);
fa40146 : full_adder port map(c30145,s30246,c30245,s40146,c40146);
fa40147 : full_adder port map(c30146,s30247,c30246,s40147,c40147);
fa40148 : full_adder port map(c30147,c10447,c30247,s40148,c40148);

--STAGE 4 GROUP 02
fa40226 : full_adder port map(s30326,c30325,c20525,s40226,c40226);
fa40228 : full_adder port map(s30328,c30327,s30428,s40228,c40228);
fa40229 : full_adder port map(s30329,c30328,s10929,s40229,c40229);
fa40230 : full_adder port map(s30330,c30329,s20630,s40230,c40230);
fa40231 : full_adder port map(s30331,c30330,s30431,s40231,c40231);
fa40232 : full_adder port map(s30332,c30331,s30432,s40232,c40232);
fa40233 : full_adder port map(s30333,c30332,s30433,s40233,c40233);
fa40234 : full_adder port map(s30334,c30333,s20634,s40234,c40234);
fa40235 : full_adder port map(s30335,c30334,s30435,s40235,c40235);
fa40236 : full_adder port map(s30336,c30335,c30435,s40236,c40236);
fa40237 : full_adder port map(s30337,c30336,c10836,s40237,c40237);
fa40238 : full_adder port map(s30338,c30337,c20537,s40238,c40238);

-----------------------------------------------------------------

--STAGE 5 -  FULL ADDERS:64 | HALF ADDERS:0
--GROUP 00
fa50007 : full_adder port map(s30007,c30006,c40006,s50007,c50007);
fa50009 : full_adder port map(s40009,c40008,c30108,s50009,c50009);
fa50011 : full_adder port map(s40011,c40010,c30110,s50011,c50011);
fa50012 : full_adder port map(s40012,c40011,c30111,s50012,c50012);
fa50013 : full_adder port map(s40013,c40012,c30112,s50013,c50013);
fa50014 : full_adder port map(s40014,c40013,c30113,s50014,c50014);
fa50015 : full_adder port map(s40015,c40014,c30114,s50015,c50015);
fa50016 : full_adder port map(s40016,c40015,s40116,s50016,c50016);
fa50017 : full_adder port map(s40017,c40016,c30116,s50017,c50017);
fa50018 : full_adder port map(s40018,c40017,s40118,s50018,c50018);
fa50019 : full_adder port map(s40019,c40018,s40119,s50019,c50019);
fa50020 : full_adder port map(s40020,c40019,s40120,s50020,c50020);
fa50021 : full_adder port map(s40021,c40020,s40121,s50021,c50021);
fa50022 : full_adder port map(s40022,c40021,s40122,s50022,c50022);
fa50023 : full_adder port map(s40023,c40022,s40123,s50023,c50023);
fa50024 : full_adder port map(s40024,c40023,s40124,s50024,c50024);
fa50025 : full_adder port map(s40025,c40024,s40125,s50025,c50025);
fa50026 : full_adder port map(s40026,c40025,s40126,s50026,c50026);
fa50027 : full_adder port map(s40027,c40026,s40127,s50027,c50027);
fa50028 : full_adder port map(s40028,c40027,s40128,s50028,c50028);
fa50029 : full_adder port map(s40029,c40028,s40129,s50029,c50029);
fa50030 : full_adder port map(s40030,c40029,s40130,s50030,c50030);
fa50031 : full_adder port map(s40031,c40030,s40131,s50031,c50031);
fa50032 : full_adder port map(s40032,c40031,s40132,s50032,c50032);
fa50033 : full_adder port map(s40033,c40032,s40133,s50033,c50033);
fa50034 : full_adder port map(s40034,c40033,s40134,s50034,c50034);
fa50035 : full_adder port map(s40035,c40034,s40135,s50035,c50035);
fa50036 : full_adder port map(s40036,c40035,s40136,s50036,c50036);
fa50037 : full_adder port map(s40037,c40036,s40137,s50037,c50037);
fa50038 : full_adder port map(s40038,c40037,s40138,s50038,c50038);
fa50039 : full_adder port map(s40039,c40038,s40139,s50039,c50039);
fa50040 : full_adder port map(s40040,c40039,s40140,s50040,c50040);
fa50041 : full_adder port map(s40041,c40040,s40141,s50041,c50041);
fa50042 : full_adder port map(s40042,c40041,s40142,s50042,c50042);
fa50043 : full_adder port map(s40043,c40042,s40143,s50043,c50043);
fa50044 : full_adder port map(s40044,c40043,s40144,s50044,c50044);
fa50045 : full_adder port map(s40045,c40044,s40145,s50045,c50045);
fa50046 : full_adder port map(s40046,c40045,s40146,s50046,c50046);
fa50047 : full_adder port map(s40047,c40046,s40147,s50047,c50047);
fa50048 : full_adder port map(s40048,c40047,s40148,s50048,c50048);
fa50049 : full_adder port map(s40049,c40048,c30148,s50049,c50049);
fa50050 : full_adder port map(s40050,c40049,c30149,s50050,c50050);
fa50051 : full_adder port map(s40051,c40050,c30150,s50051,c50051);
fa50052 : full_adder port map(s40052,c40051,c30151,s50052,c50052);
fa50053 : full_adder port map(s40053,c40052,c30152,s50053,c50053);
fa50054 : full_adder port map(s40054,c40053,c30153,s50054,c50054);
fa50056 : full_adder port map(s40056,c40055,c30155,s50056,c50056);
fa50059 : full_adder port map(s30059,c30058,c40058,s50059,c50059);

--STAGE 5 GROUP 01
fa50123 : full_adder port map(c40122,c20422,c30322,s50123,c50123);
fa50125 : full_adder port map(c40124,s30325,c30324,s50125,c50125);
fa50127 : full_adder port map(c40126,s30327,c30326,s50127,c50127);
fa50129 : full_adder port map(c40128,s40229,c40228,s50129,c50129);
fa50130 : full_adder port map(c40129,s40230,c40229,s50130,c50130);
fa50131 : full_adder port map(c40130,s40231,c40230,s50131,c50131);
fa50132 : full_adder port map(c40131,s40232,c40231,s50132,c50132);
fa50133 : full_adder port map(c40132,s40233,c40232,s50133,c50133);
fa50134 : full_adder port map(c40133,s40234,c40233,s50134,c50134);
fa50135 : full_adder port map(c40134,s40235,c40234,s50135,c50135);
fa50136 : full_adder port map(c40135,s40236,c40235,s50136,c50136);
fa50137 : full_adder port map(c40136,s40237,c40236,s50137,c50137);
fa50138 : full_adder port map(c40137,s40238,c40237,s50138,c50138);
fa50139 : full_adder port map(c40138,s30339,c30338,s50139,c50139);
fa50140 : full_adder port map(c40139,s30340,c30339,s50140,c50140);
fa50141 : full_adder port map(c40140,c20440,c30340,s50141,c50141);

-----------------------------------------------------------------

--STAGE 6 -  FULL ADDERS:40 | HALF ADDERS:0
--GROUP 00
fa60010 : full_adder port map(s40010,c40009,c50009,s60010,c60010);
fa60013 : full_adder port map(s50013,c50012,p(416),s60013,c60013);
fa60015 : full_adder port map(s50015,c50014,s30215,s60015,c60015);
fa60017 : full_adder port map(s50017,c50016,s30217,s60017,c60017);
fa60019 : full_adder port map(s50019,c50018,c40118,s60019,c60019);
fa60020 : full_adder port map(s50020,c50019,c40119,s60020,c60020);
fa60021 : full_adder port map(s50021,c50020,c40120,s60021,c60021);
fa60022 : full_adder port map(s50022,c50021,c40121,s60022,c60022);
fa60023 : full_adder port map(s50023,c50022,s50123,s60023,c60023);
fa60024 : full_adder port map(s50024,c50023,c40123,s60024,c60024);
fa60025 : full_adder port map(s50025,c50024,s50125,s60025,c60025);
fa60026 : full_adder port map(s50026,c50025,c40125,s60026,c60026);
fa60027 : full_adder port map(s50027,c50026,s50127,s60027,c60027);
fa60028 : full_adder port map(s50028,c50027,c40127,s60028,c60028);
fa60029 : full_adder port map(s50029,c50028,s50129,s60029,c60029);
fa60030 : full_adder port map(s50030,c50029,s50130,s60030,c60030);
fa60031 : full_adder port map(s50031,c50030,s50131,s60031,c60031);
fa60032 : full_adder port map(s50032,c50031,s50132,s60032,c60032);
fa60033 : full_adder port map(s50033,c50032,s50133,s60033,c60033);
fa60034 : full_adder port map(s50034,c50033,s50134,s60034,c60034);
fa60035 : full_adder port map(s50035,c50034,s50135,s60035,c60035);
fa60036 : full_adder port map(s50036,c50035,s50136,s60036,c60036);
fa60037 : full_adder port map(s50037,c50036,s50137,s60037,c60037);
fa60038 : full_adder port map(s50038,c50037,s50138,s60038,c60038);
fa60039 : full_adder port map(s50039,c50038,s50139,s60039,c60039);
fa60040 : full_adder port map(s50040,c50039,s50140,s60040,c60040);
fa60041 : full_adder port map(s50041,c50040,s50141,s60041,c60041);
fa60042 : full_adder port map(s50042,c50041,c40141,s60042,c60042);
fa60043 : full_adder port map(s50043,c50042,c40142,s60043,c60043);
fa60044 : full_adder port map(s50044,c50043,c40143,s60044,c60044);
fa60045 : full_adder port map(s50045,c50044,c40144,s60045,c60045);
fa60046 : full_adder port map(s50046,c50045,c40145,s60046,c60046);
fa60047 : full_adder port map(s50047,c50046,c40146,s60047,c60047);
fa60048 : full_adder port map(s50048,c50047,c40147,s60048,c60048);
fa60049 : full_adder port map(s50049,c50048,s30249,s60049,c60049);
fa60050 : full_adder port map(s50050,c50049,c30249,s60050,c60050);
fa60051 : full_adder port map(s50051,c50050,c20250,s60051,c60051);
fa60055 : full_adder port map(s40055,c40054,c50054,s60055,c60055);
fa60057 : full_adder port map(s40057,c40056,c50056,s60057,c60057);
fa60060 : full_adder port map(s30060,c30059,c50059,s60060,c60060);

-----------------------------------------------------------------

--STAGE 7 -  FULL ADDERS:28 | HALF ADDERS:0
--GROUP 00
fa70014 : full_adder port map(s50014,c50013,c60013,s70014,c70014);
fa70016 : full_adder port map(s50016,c50015,c60015,s70016,c70016);
fa70018 : full_adder port map(s50018,c50017,c60017,s70018,c70018);
fa70022 : full_adder port map(s60022,c60021,s30322,s70022,c70022);
fa70024 : full_adder port map(s60024,c60023,s30324,s70024,c70024);
fa70026 : full_adder port map(s60026,c60025,s40226,s70026,c70026);
fa70027 : full_adder port map(s60027,c60026,c40226,s70027,c70027);
fa70028 : full_adder port map(s60028,c60027,s40228,s70028,c70028);
fa70029 : full_adder port map(s60029,c60028,c30428,s70029,c70029);
fa70030 : full_adder port map(s60030,c60029,c50129,s70030,c70030);
fa70031 : full_adder port map(s60031,c60030,c50130,s70031,c70031);
fa70032 : full_adder port map(s60032,c60031,c50131,s70032,c70032);
fa70033 : full_adder port map(s60033,c60032,c50132,s70033,c70033);
fa70034 : full_adder port map(s60034,c60033,c50133,s70034,c70034);
fa70035 : full_adder port map(s60035,c60034,c50134,s70035,c70035);
fa70036 : full_adder port map(s60036,c60035,c50135,s70036,c70036);
fa70037 : full_adder port map(s60037,c60036,c50136,s70037,c70037);
fa70038 : full_adder port map(s60038,c60037,c50137,s70038,c70038);
fa70039 : full_adder port map(s60039,c60038,c50138,s70039,c70039);
fa70040 : full_adder port map(s60040,c60039,c50139,s70040,c70040);
fa70041 : full_adder port map(s60041,c60040,c50140,s70041,c70041);
fa70042 : full_adder port map(s60042,c60041,s30342,s70042,c70042);
fa70043 : full_adder port map(s60043,c60042,c30342,s70043,c70043);
fa70044 : full_adder port map(s60044,c60043,c20443,s70044,c70044);
fa70049 : full_adder port map(s60049,c60048,c40148,s70049,c70049);
fa70052 : full_adder port map(s50052,c50051,c60051,s70052,c70052);
fa70058 : full_adder port map(s40058,c40057,c60057,s70058,c70058);
fa70061 : full_adder port map(s20061,c30060,c60060,s70061,c70061);

-----------------------------------------------------------------

--STAGE 8 -  FULL ADDERS:14 | HALF ADDERS:21
--GROUP 00
fa80017 : full_adder port map(s60017,c40116,c70016,s80017,c80017);
fa80019 : full_adder port map(s60019,p(608),c70018,s80019,c80019);
ha80020 : half_adder port map(s60020,c60019,s80020,c80020);
ha80021 : half_adder port map(s60021,c60020,s80021,c80021);
fa80023 : full_adder port map(s60023,c60022,c70022,s80023,c80023);
ha80024 : half_adder port map(s70024,c50123,s80024,c80024);
fa80025 : full_adder port map(s60025,c60024,c70024,s80025,c80025);
ha80026 : half_adder port map(s70026,c50125,s80026,c80026);
ha80027 : half_adder port map(s70027,c70026,s80027,c80027);
fa80028 : full_adder port map(s70028,c70027,c50127,s80028,c80028);
ha80029 : half_adder port map(s70029,c70028,s80029,c80029);
ha80030 : half_adder port map(s70030,c70029,s80030,c80030);
ha80031 : half_adder port map(s70031,c70030,s80031,c80031);
fa80032 : full_adder port map(s70032,c70031,c30431,s80032,c80032);
fa80033 : full_adder port map(s70033,c70032,c30432,s80033,c80033);
fa80034 : full_adder port map(s70034,c70033,c30433,s80034,c80034);
ha80035 : half_adder port map(s70035,c70034,s80035,c80035);
ha80036 : half_adder port map(s70036,c70035,s80036,c80036);
ha80037 : half_adder port map(s70037,c70036,s80037,c80037);
ha80038 : half_adder port map(s70038,c70037,s80038,c80038);
fa80039 : full_adder port map(s70039,c70038,c40238,s80039,c80039);
ha80040 : half_adder port map(s70040,c70039,s80040,c80040);
ha80041 : half_adder port map(s70041,c70040,s80041,c80041);
fa80042 : full_adder port map(s70042,c70041,c50141,s80042,c80042);
ha80043 : half_adder port map(s70043,c70042,s80043,c80043);
ha80044 : half_adder port map(s70044,c70043,s80044,c80044);
fa80045 : full_adder port map(s60045,c60044,c70044,s80045,c80045);
ha80046 : half_adder port map(s60046,c60045,s80046,c80046);
ha80047 : half_adder port map(s60047,c60046,s80047,c80047);
ha80048 : half_adder port map(s60048,c60047,s80048,c80048);
fa80050 : full_adder port map(s60050,c60049,c70049,s80050,c80050);
ha80051 : half_adder port map(s60051,c60050,s80051,c80051);
fa80053 : full_adder port map(s50053,c50052,c70052,s80053,c80053);
ha80054 : half_adder port map(s50054,c50053,s80054,c80054);
fa80062 : full_adder port map(p(1023),c20061,c70061,s80062,c80062);